module DiffBridge(
  input        clock,
  input [ 7:0] coreid,

  input [ 7:0] index_0,
  input        Instrvalid_0,
  input [63:0] the_pc_0,
  input [31:0] instr_0,
  input        skip_0,
  input        is_TLBFILL_0,
  input [ 4:0] TLBFILL_index_0,
  input        is_CNTinst_0,
  input [63:0] timer_64_value_0,
  input        wen_0,
  input [ 7:0] wdest_0,
  input [63:0] wdata_0,
  input        csr_rstat_0,
  input [31:0] csr_data_0,

  input [ 7:0] index_1,
  input        Instrvalid_1,
  input [63:0] the_pc_1,
  input [31:0] instr_1,
  input        skip_1,
  input        is_TLBFILL_1,
  input [ 4:0] TLBFILL_index_1,
  input        is_CNTinst_1,
  input [63:0] timer_64_value_1,
  input        wen_1,
  input [ 7:0] wdest_1,
  input [63:0] wdata_1,
  input        csr_rstat_1,
  input [31:0] csr_data_1,

  input [ 7:0] index_2,
  input        Instrvalid_2,
  input [63:0] the_pc_2,
  input [31:0] instr_2,
  input        skip_2,
  input        is_TLBFILL_2,
  input [ 4:0] TLBFILL_index_2,
  input        is_CNTinst_2,
  input [63:0] timer_64_value_2,
  input        wen_2,
  input [ 7:0] wdest_2,
  input [63:0] wdata_2,
  input        csr_rstat_2,
  input [31:0] csr_data_2,
  
  input [ 7:0] index_3,
  input        Instrvalid_3,
  input [63:0] the_pc_3,
  input [31:0] instr_3,
  input        skip_3,
  input        is_TLBFILL_3,
  input [ 4:0] TLBFILL_index_3,
  input        is_CNTinst_3,
  input [63:0] timer_64_value_3,
  input        wen_3,
  input [ 7:0] wdest_3,
  input [63:0] wdata_3,
  input        csr_rstat_3,
  input [31:0] csr_data_3,

  input [ 7:0] storeIndex,
  input [ 7:0] storeValid,
  input [63:0] storePaddr,
  input [63:0] storeVaddr,
  input [63:0] storeData,

  input [63:0] REG_0,
  input [63:0] REG_1,
  input [63:0] REG_2,
  input [63:0] REG_3,
  input [63:0] REG_4,
  input [63:0] REG_5,
  input [63:0] REG_6,
  input [63:0] REG_7,
  input [63:0] REG_8,
  input [63:0] REG_9,
  input [63:0] REG_10,
  input [63:0] REG_11,
  input [63:0] REG_12,
  input [63:0] REG_13,
  input [63:0] REG_14,
  input [63:0] REG_15,
  input [63:0] REG_16,
  input [63:0] REG_17,
  input [63:0] REG_18,
  input [63:0] REG_19,
  input [63:0] REG_20,
  input [63:0] REG_21,
  input [63:0] REG_22,
  input [63:0] REG_23,
  input [63:0] REG_24,
  input [63:0] REG_25,
  input [63:0] REG_26,
  input [63:0] REG_27,
  input [63:0] REG_28,
  input [63:0] REG_29,
  input [63:0] REG_30,
  input [63:0] REG_31
);

DifftestInstrCommit DifftestInstrCommit_0(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .index              (index_0        ),
  .valid              (Instrvalid_0   ),
  .pc                 (the_pc_0       ),
  .instr              (instr_0        ),
  .skip               (skip_0         ),
  .is_TLBFILL         (is_TLBFILL_0   ),
  .TLBFILL_index      (TLBFILL_index_0),
  .is_CNTinst         (is_CNTinst_0   ),
  .timer_64_value     (timer_64_value_0),
  .wen                (wen_0          ),
  .wdest              (wdest_0        ),
  .wdata              (wdata_0        ),
  .csr_rstat          (csr_rstat_0    ),
  .csr_data           (csr_data_0     )
);

DifftestInstrCommit DifftestInstrCommit_1(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .index              (index_1        ),
  .valid              (Instrvalid_1   ),
  .pc                 (the_pc_1       ),
  .instr              (instr_1        ),
  .skip               (skip_1         ),
  .is_TLBFILL         (is_TLBFILL_1   ),
  .TLBFILL_index      (TLBFILL_index_1),
  .is_CNTinst         (is_CNTinst_1   ),
  .timer_64_value     (timer_64_value_1),
  .wen                (wen_1          ),
  .wdest              (wdest_1        ),
  .wdata              (wdata_1        ),
  .csr_rstat          (csr_rstat_1    ),
  .csr_data           (csr_data_1     )
);

DifftestInstrCommit DifftestInstrCommit_2(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .index              (index_2        ),
  .valid              (Instrvalid_2   ),
  .pc                 (the_pc_2       ),
  .instr              (instr_2        ),
  .skip               (skip_2         ),
  .is_TLBFILL         (is_TLBFILL_2   ),
  .TLBFILL_index      (TLBFILL_index_2),
  .is_CNTinst         (is_CNTinst_2   ),
  .timer_64_value     (timer_64_value_2),
  .wen                (wen_2          ),
  .wdest              (wdest_2        ),
  .wdata              (wdata_2        ),
  .csr_rstat          (csr_rstat_2    ),
  .csr_data           (csr_data_2     )
);

DifftestInstrCommit DifftestInstrCommit_3(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .index              (index_3        ),
  .valid              (Instrvalid_3   ),
  .pc                 (the_pc_3       ),
  .instr              (instr_3        ),
  .skip               (skip_3         ),
  .is_TLBFILL         (is_TLBFILL_3   ),
  .TLBFILL_index      (TLBFILL_index_3),
  .is_CNTinst         (is_CNTinst_3   ),
  .timer_64_value     (timer_64_value_3),
  .wen                (wen_3          ),
  .wdest              (wdest_3        ),
  .wdata              (wdata_3        ),
  .csr_rstat          (csr_rstat_3    ),
  .csr_data           (csr_data_3     )
);

DifftestStoreEvent DifftestStoreEvent_1(
  .clock              (clock          ),
  .coreid             (0              ),
  .index              (storeIndex   ),
  .valid              (storeValid   ),
  .storePAddr         (storePaddr   ),
  .storeVAddr         (storeVaddr   ),
  .storeData          (storeData    )
);

DifftestGRegState DifftestGRegState_0(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .gpr_0              (REG_0          ),
  .gpr_1              (REG_1          ),
  .gpr_2              (REG_2          ),
  .gpr_3              (REG_3          ),
  .gpr_4              (REG_4          ),
  .gpr_5              (REG_5          ),
  .gpr_6              (REG_6          ),
  .gpr_7              (REG_7          ),
  .gpr_8              (REG_8          ),
  .gpr_9              (REG_9          ),
  .gpr_10             (REG_10         ),
  .gpr_11             (REG_11         ),
  .gpr_12             (REG_12         ),
  .gpr_13             (REG_13         ),
  .gpr_14             (REG_14         ),
  .gpr_15             (REG_15         ),
  .gpr_16             (REG_16         ),
  .gpr_17             (REG_17         ),
  .gpr_18             (REG_18         ),
  .gpr_19             (REG_19         ),
  .gpr_20             (REG_20         ),
  .gpr_21             (REG_21         ),
  .gpr_22             (REG_22         ),
  .gpr_23             (REG_23         ),
  .gpr_24             (REG_24         ),
  .gpr_25             (REG_25         ),
  .gpr_26             (REG_26         ),
  .gpr_27             (REG_27         ),
  .gpr_28             (REG_28         ),
  .gpr_29             (REG_29         ),
  .gpr_30             (REG_30         ),
  .gpr_31             (REG_31         )
);

endmodule
