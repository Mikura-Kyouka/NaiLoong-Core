module DiffBridge(
  input        clock,
  input [ 7:0] coreid,

  input [ 7:0] index_0,
  input        Instrvalid_0,
  input [63:0] the_pc_0,
  input [31:0] instr_0,
  input        skip_0,
  input        is_TLBFILL_0,
  input [ 4:0] TLBFILL_index_0,
  input        is_CNTinst_0,
  input [63:0] timer_64_value_0,
  input        wen_0,
  input [ 7:0] wdest_0,
  input [63:0] wdata_0,
  input        csr_rstat_0,
  input [31:0] csr_data_0,

  input [ 7:0] index_1,
  input        Instrvalid_1,
  input [63:0] the_pc_1,
  input [31:0] instr_1,
  input        skip_1,
  input        is_TLBFILL_1,
  input [ 4:0] TLBFILL_index_1,
  input        is_CNTinst_1,
  input [63:0] timer_64_value_1,
  input        wen_1,
  input [ 7:0] wdest_1,
  input [63:0] wdata_1,
  input        csr_rstat_1,
  input [31:0] csr_data_1,

  input [ 7:0] index_2,
  input        Instrvalid_2,
  input [63:0] the_pc_2,
  input [31:0] instr_2,
  input        skip_2,
  input        is_TLBFILL_2,
  input [ 4:0] TLBFILL_index_2,
  input        is_CNTinst_2,
  input [63:0] timer_64_value_2,
  input        wen_2,
  input [ 7:0] wdest_2,
  input [63:0] wdata_2,
  input        csr_rstat_2,
  input [31:0] csr_data_2,

  input        excp_valid,
  input        eret,
  input [10:0] intrNo,
  input [ 5:0] cause,
  input [31:0] exceptionPC,
  input [31:0] exceptionInst,

  input [ 7:0] storeIndex,
  input [ 7:0] storeValid,
  input [63:0] storePaddr,
  input [63:0] storeVaddr,
  input [63:0] storeData,

  input [ 7:0] loadIndex,
  input [ 7:0] loadValid,
  input [63:0] loadPaddr,
  input [63:0] loadVaddr,

  input [63:0] REG_0,
  input [63:0] REG_1,
  input [63:0] REG_2,
  input [63:0] REG_3,
  input [63:0] REG_4,
  input [63:0] REG_5,
  input [63:0] REG_6,
  input [63:0] REG_7,
  input [63:0] REG_8,
  input [63:0] REG_9,
  input [63:0] REG_10,
  input [63:0] REG_11,
  input [63:0] REG_12,
  input [63:0] REG_13,
  input [63:0] REG_14,
  input [63:0] REG_15,
  input [63:0] REG_16,
  input [63:0] REG_17,
  input [63:0] REG_18,
  input [63:0] REG_19,
  input [63:0] REG_20,
  input [63:0] REG_21,
  input [63:0] REG_22,
  input [63:0] REG_23,
  input [63:0] REG_24,
  input [63:0] REG_25,
  input [63:0] REG_26,
  input [63:0] REG_27,
  input [63:0] REG_28,
  input [63:0] REG_29,
  input [63:0] REG_30,
  input [63:0] REG_31,

  input [63:0] CSR_0,
  input [63:0] CSR_1,
  input [63:0] CSR_2,
  input [63:0] CSR_3,
  input [63:0] CSR_4,
  input [63:0] CSR_5,
  input [63:0] CSR_6,
  input [63:0] CSR_7,
  input [63:0] CSR_8,
  input [63:0] CSR_9,
  input [63:0] CSR_10,
  input [63:0] CSR_11,
  input [63:0] CSR_12,
  input [63:0] CSR_13,
  input [63:0] CSR_14,
  input [63:0] CSR_15,
  input [63:0] CSR_16,
  input [63:0] CSR_17,
  input [63:0] CSR_18,
  input [63:0] CSR_19,
  input [63:0] CSR_20,
  input [63:0] CSR_21,
  input [63:0] CSR_22,
  input [63:0] CSR_23,
  input [63:0] CSR_24,
  input [63:0] CSR_25,
  input [63:0] CSR_26
);

DifftestExcpEvent DifftestExcpEvent(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .excp_valid         (excp_valid     ),
  .eret               (eret           ),
  .intrNo             (intrNo         ),
  .cause              (cause          ),
  .exceptionPC        (exceptionPC    ),
  .exceptionInst      (exceptionInst  )
);

DifftestInstrCommit DifftestInstrCommit_0(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .index              (index_0        ),
  .valid              (Instrvalid_0   ),
  .pc                 (the_pc_0       ),
  .instr              (instr_0        ),
  .skip               (skip_0         ),
  .is_TLBFILL         (is_TLBFILL_0   ),
  .TLBFILL_index      (TLBFILL_index_0),
  .is_CNTinst         (is_CNTinst_0   ),
  .timer_64_value     (timer_64_value_0),
  .wen                (wen_0          ),
  .wdest              (wdest_0        ),
  .wdata              (wdata_0        ),
  .csr_rstat          (csr_rstat_0    ),
  .csr_data           (csr_data_0     )
);

DifftestInstrCommit DifftestInstrCommit_1(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .index              (index_1        ),
  .valid              (Instrvalid_1   ),
  .pc                 (the_pc_1       ),
  .instr              (instr_1        ),
  .skip               (skip_1         ),
  .is_TLBFILL         (is_TLBFILL_1   ),
  .TLBFILL_index      (TLBFILL_index_1),
  .is_CNTinst         (is_CNTinst_1   ),
  .timer_64_value     (timer_64_value_1),
  .wen                (wen_1          ),
  .wdest              (wdest_1        ),
  .wdata              (wdata_1        ),
  .csr_rstat          (csr_rstat_1    ),
  .csr_data           (csr_data_1     )
);

// DifftestInstrCommit DifftestInstrCommit_2(
//   .clock              (clock          ),
//   .coreid             (coreid         ),
//   .index              (index_2        ),
//   .valid              (Instrvalid_2   ),
//   .pc                 (the_pc_2       ),
//   .instr              (instr_2        ),
//   .skip               (skip_2         ),
//   .is_TLBFILL         (is_TLBFILL_2   ),
//   .TLBFILL_index      (TLBFILL_index_2),
//   .is_CNTinst         (is_CNTinst_2   ),
//   .timer_64_value     (timer_64_value_2),
//   .wen                (wen_2          ),
//   .wdest              (wdest_2        ),
//   .wdata              (wdata_2        ),
//   .csr_rstat          (csr_rstat_2    ),
//   .csr_data           (csr_data_2     )
// );

DifftestStoreEvent DifftestStoreEvent_1(
  .clock              (clock          ),
  .coreid             (0              ),
  .index              (storeIndex   ),
  .valid              (storeValid   ),
  .storePAddr         (storePaddr   ),
  .storeVAddr         (storeVaddr   ),
  .storeData          (storeData    )
);

DifftestLoadEvent DifftestLoadEvent_1(
  .clock              (clock          ),
  .coreid             (0              ),
  .index              (loadIndex      ),
  .valid              (loadValid      ),
  .paddr              (loadPaddr      ),
  .vaddr              (loadVaddr      )
);

DifftestGRegState DifftestGRegState_0(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .gpr_0              (REG_0          ),
  .gpr_1              (REG_1          ),
  .gpr_2              (REG_2          ),
  .gpr_3              (REG_3          ),
  .gpr_4              (REG_4          ),
  .gpr_5              (REG_5          ),
  .gpr_6              (REG_6          ),
  .gpr_7              (REG_7          ),
  .gpr_8              (REG_8          ),
  .gpr_9              (REG_9          ),
  .gpr_10             (REG_10         ),
  .gpr_11             (REG_11         ),
  .gpr_12             (REG_12         ),
  .gpr_13             (REG_13         ),
  .gpr_14             (REG_14         ),
  .gpr_15             (REG_15         ),
  .gpr_16             (REG_16         ),
  .gpr_17             (REG_17         ),
  .gpr_18             (REG_18         ),
  .gpr_19             (REG_19         ),
  .gpr_20             (REG_20         ),
  .gpr_21             (REG_21         ),
  .gpr_22             (REG_22         ),
  .gpr_23             (REG_23         ),
  .gpr_24             (REG_24         ),
  .gpr_25             (REG_25         ),
  .gpr_26             (REG_26         ),
  .gpr_27             (REG_27         ),
  .gpr_28             (REG_28         ),
  .gpr_29             (REG_29         ),
  .gpr_30             (REG_30         ),
  .gpr_31             (REG_31         )
);

DifftestCSRRegState DifftestCSRRegState_0(
  .clock              (clock          ),
  .coreid             (coreid         ),
  .crmd               (CSR_0          ),
  .prmd               (CSR_1          ),
  .euen               (CSR_2          ),
  .ecfg               (CSR_3          ),
  .estat              (CSR_4          ),
  .era                (CSR_5          ),
  .badv               (CSR_6          ),
  .eentry             (CSR_7          ),
  .tlbidx             (CSR_8          ),
  .tlbehi             (CSR_9          ),
  .tlbelo0            (CSR_10         ),
  .tlbelo1            (CSR_11         ),
  .asid               (CSR_12         ),
  .pgdl               (CSR_13         ),
  .pgdh               (CSR_14         ),
  .save0              (CSR_15         ),
  .save1              (CSR_16         ),
  .save2              (CSR_17         ),
  .save3              (CSR_18         ),
  .tid                (CSR_19         ),
  .tcfg               (CSR_20         ),
  .tval               (CSR_21         ),
  .ticlr              (CSR_22         ),
  .llbctl             (CSR_23         ),
  .tlbrentry          (CSR_24         ),
  .dmw0               (CSR_25         ),
  .dmw1               (CSR_26         )
);

endmodule
